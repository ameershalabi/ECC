--------------------------------------------------------------------------------
-- Title       : Hamming Package
-- Project     : ECC 
--------------------------------------------------------------------------------
-- File        : hamming_pkg.vhd
-- Author      : Ameer Shalabi <ameershalabi94@gmail.com>
-- Company     : User Company Name
-- Created     : Sat Oct 26 11:03:09 2024
-- Last update : Sun Nov 10 11:41:04 2024
-- Platform    : -
-- Standard    : <VHDL-2008 | VHDL-2002 | VHDL-1993 | VHDL-1987>
--------------------------------------------------------------------------------
-- Copyright (c) 2024 User Company Name
-------------------------------------------------------------------------------
-- Description: 
--------------------------------------------------------------------------------
-- Revisions:  Revisions and documentation are controlled by
-- the revision control system (RCS).  The RCS should be consulted
-- on revision history.
-------------------------------------------------------------------------------
library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package hamming_pkg is

  constant parity_0_loc_placement : std_logic_vector(523 downto 0) :=
    x"15555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555";
  ----00010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010
  ----10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101
  ----01010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010
  ----10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101
  constant parity_1_loc_placement : std_logic_vector(523 downto 0) :=
    x"26666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666";
  ----00100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011
  ----00110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001
  ----10011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100
  ----11001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110
  constant parity_3_loc_placement : std_logic_vector(523 downto 0) :=
    x"07878787878787878787878787878787878787878787878787878787878787878787878787878787878787878787878787878787878787878787878787878787878";
  ----00000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100
  ----00111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001
  ----11100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111
  ----00001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000
  constant parity_7_loc_placement : std_logic_vector(523 downto 0) :=
    x"3807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f807f80";
  ----00111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111
  ----11000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110
  ----00000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000
  ----00001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000
  constant parity_15_loc_placement : std_logic_vector(523 downto 0) :=
    x"0007fff80007fff80007fff80007fff80007fff80007fff80007fff80007fff80007fff80007fff80007fff80007fff80007fff80007fff80007fff80007fff8000";
  ----00000000000001111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000
  ----00000000001111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000
  ----00000001111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000
  ----00001111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000
  constant parity_31_loc_placement : std_logic_vector(523 downto 0) :=
    x"0007fffffff800000007fffffff800000007fffffff800000007fffffff800000007fffffff800000007fffffff800000007fffffff800000007fffffff80000000";
  ----00000000000001111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000
  ----00000000001111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000
  ----00000001111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000
  ----00001111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000
  constant parity_63_loc_placement : std_logic_vector(523 downto 0) :=
    x"0007fffffffffffffff80000000000000007fffffffffffffff80000000000000007fffffffffffffff80000000000000007fffffffffffffff8000000000000000";
  ----00000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000
  ----00000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000
  ----00000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000
  ----00001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000
  constant parity_127_loc_placement : std_logic_vector(523 downto 0) :=
    x"0007fffffffffffffffffffffffffffffff800000000000000000000000000000007fffffffffffffffffffffffffffffff80000000000000000000000000000000";
  ----00000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
  ----11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
  ----00000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
  ----11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
  constant parity_255_loc_placement : std_logic_vector(523 downto 0) :=
    x"0007fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8000000000000000000000000000000000000000000000000000000000000000";
  ----00000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
  ----11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
  ----11111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
  ----00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000

  constant parity_511_loc_placement : std_logic_vector(523 downto 0) :=
    x"3ff80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  ----00111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
  ----00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
  ----00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
  ----00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000

  function num_parity_bits (data_w : integer) return integer;
  function generate_xor_tree_logic (data : std_logic_vector) return std_logic;
  function count_1s (vector        : std_logic_vector) return natural;

  -- arr to hold xor results of tree_depth x w_position_vector
  type xor_tree_t is array (integer range <>,
      integer range <>) of std_logic;

end package hamming_pkg;

-- Package Body Section
package body hamming_pkg is

  function num_parity_bits (data_w : integer) return integer is
    variable n_parity : integer := 0;
  begin
    get_number_of_parity : while (2**n_parity < data_w + n_parity + 1) loop
      n_parity := n_parity +1;
    end loop get_number_of_parity;
    return n_parity;
  end function num_parity_bits;

  function count_1s (vector : std_logic_vector) return natural is
    variable count : natural := 0;
  begin
    loop_over_data : for i in 0 to vector'length-1 loop
      if vector(i) = '1' then
        count := count+1;
      end if;
    end loop loop_over_data;
    return count;
  end function count_1s;

  function generate_xor_tree_logic (
      data : std_logic_vector
    )
    return std_logic is
    variable depth_xor_tree : positive := positive(ceil(log2(real(data'length))));
    variable xor_tree       : xor_tree_t(0 to depth_xor_tree,0 to data'length-1);
    variable nodes_per_depth : integer range 0 to data'length-1;
  begin
    max_depth_data_loop : for b in 0 to data'length-1 loop
      xor_tree(depth_xor_tree,b)  := data(b);
    end loop max_depth_data_loop;

    dpeth_loop : for depth in depth_xor_tree-1 downto 0 loop
      nodes_per_depth:= 2**depth;
      nodes_loop : for node in 0 to nodes_per_depth-1 loop
        xor_tree(depth,node) :=  xor_tree(depth+1,node*2) xor  xor_tree(depth+1,node*2 +1);
      end loop nodes_loop;
    end loop dpeth_loop;
  return xor_tree(0,0);
  end function generate_xor_tree_logic;

end package body hamming_pkg;